module twiddle_factor_rom (input logic [10:0] addr_t,
									output logic [31:0] twiddle);
	parameter ADDR_WIDTH = 11;
   parameter DATA_WIDTH =  32;
	logic [ADDR_WIDTH-1:0] addr_reg;

	parameter [0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM0 = {
		32'b01111111111111110000000000000000,
		32'b01111111111111110000000001100100,
		32'b01111111111111110000000011001001,
		32'b01111111111111100000000100101101,
		32'b01111111111111010000000110010010,
		32'b01111111111111000000000111110110,
		32'b01111111111110100000001001011011,
		32'b01111111111110000000001010111111,
		32'b01111111111101100000001100100100,
		32'b01111111111100110000001110001000,
		32'b01111111111100000000001111101101,
		32'b01111111111011010000010001010001,
		32'b01111111111010010000010010110110,
		32'b01111111111001010000010100011010,
		32'b01111111111000010000010101111111,
		32'b01111111110111010000010111100011,
		32'b01111111110110000000011001000111,
		32'b01111111110100110000011010101100,
		32'b01111111110011100000011100010000,
		32'b01111111110010000000011101110101,
		32'b01111111110000100000011111011001,
		32'b01111111101111000000100000111101,
		32'b01111111101101010000100010100010,
		32'b01111111101011100000100100000110,
		32'b01111111101001110000100101101010,
		32'b01111111100111110000100111001110,
		32'b01111111100101110000101000110011,
		32'b01111111100011110000101010010111,
		32'b01111111100001110000101011111011,
		32'b01111111011111100000101101011111,
		32'b01111111011101010000101111000011,
		32'b01111111011010110000110000100111,
		32'b01111111011000100000110010001011,
		32'b01111111010110000000110011101111,
		32'b01111111010011010000110101010011,
		32'b01111111010000110000110110110111,
		32'b01111111001110000000111000011011,
		32'b01111111001011010000111001111111,
		32'b01111111001000010000111011100011,
		32'b01111111000101010000111101000111,
		32'b01111111000010010000111110101011,
		32'b01111110111111010001000000001110,
		32'b01111110111100000001000001110010,
		32'b01111110111000110001000011010110,
		32'b01111110110101010001000100111001,
		32'b01111110110010000001000110011101,
		32'b01111110101110100001001000000001,
		32'b01111110101010110001001001100100,
		32'b01111110100111010001001011001000,
		32'b01111110100011100001001100101011,
		32'b01111110011111110001001110001110,
		32'b01111110011011110001001111110010,
		32'b01111110010111110001010001010101,
		32'b01111110010011110001010010111000,
		32'b01111110001111110001010100011011,
		32'b01111110001011100001010101111111,
		32'b01111110000111010001010111100010,
		32'b01111110000011000001011001000101,
		32'b01111101111110100001011010101000,
		32'b01111101111010000001011100001010,
		32'b01111101110101100001011101101101,
		32'b01111101110000110001011111010000,
		32'b01111101101100000001100000110011,
		32'b01111101100111010001100010010110,
		32'b01111101100010100001100011111000,
		32'b01111101011101100001100101011011,
		32'b01111101011000100001100110111101,
		32'b01111101010011100001101000100000,
		32'b01111101001110010001101010000010,
		32'b01111101001001000001101011100100,
		32'b01111101000011110001101101000111,
		32'b01111100111110010001101110101001,
		32'b01111100111000110001110000001011,
		32'b01111100110011010001110001101101,
		32'b01111100101101110001110011001111,
		32'b01111100101000000001110100110001,
		32'b01111100100010010001110110010011,
		32'b01111100011100010001110111110101,
		32'b01111100010110100001111001010110,
		32'b01111100010000100001111010111000,
		32'b01111100001010010001111100011001,
		32'b01111100000100010001111101111011,
		32'b01111011111110000001111111011100,
		32'b01111011110111110010000000111110,
		32'b01111011110001010010000010011111,
		32'b01111011101011000010000100000000,
		32'b01111011100100100010000101100001,
		32'b01111011011101110010000111000010,
		32'b01111011010111010010001000100011,
		32'b01111011010000100010001010000100,
		32'b01111011001001100010001011100101,
		32'b01111011000010110010001101000101,
		32'b01111010111011110010001110100110,
		32'b01111010110100110010010000000111,
		32'b01111010101101100010010001100111,
		32'b01111010100110100010010011000111,
		32'b01111010011111010010010100101000,
		32'b01111010010111110010010110001000,
		32'b01111010010000100010010111101000,
		32'b01111010001001000010011001001000,
		32'b01111010000001010010011010101000,
		32'b01111001111001110010011100000111,
		32'b01111001110010000010011101100111,
		32'b01111001101010010010011111000111,
		32'b01111001100010100010100000100110,
		32'b01111001011010100010100010000110,
		32'b01111001010010100010100011100101,
		32'b01111001001010100010100101000100,
		32'b01111001000010010010100110100011,
		32'b01111000111010000010101000000010,
		32'b01111000110001110010101001100001,
		32'b01111000101001100010101011000000,
		32'b01111000100001000010101100011111,
		32'b01111000011000100010101101111101,
		32'b01111000010000000010101111011100,
		32'b01111000000111010010110000111010,
		32'b01110111111110100010110010011000,
		32'b01110111110101110010110011110111,
		32'b01110111101101000010110101010101,
		32'b01110111100100000010110110110011,
		32'b01110111011011000010111000010001,
		32'b01110111010001110010111001101110,
		32'b01110111001000110010111011001100,
		32'b01110110111111100010111100101001,
		32'b01110110110110010010111110000111,
		32'b01110110101100110010111111100100,
		32'b01110110100011100011000001000001,
		32'b01110110011010000011000010011110,
		32'b01110110010000010011000011111011,
		32'b01110110000110110011000101011000,
		32'b01110101111101000011000110110101,
		32'b01110101110011000011001000010001,
		32'b01110101101001010011001001101110,
		32'b01110101011111010011001011001010,
		32'b01110101010101010011001100100110,
		32'b01110101001011010011001110000010,
		32'b01110101000001000011001111011110,
		32'b01110100110110110011010000111010,
		32'b01110100101100100011010010010110,
		32'b01110100100010010011010011110010,
		32'b01110100010111110011010101001101,
		32'b01110100001101010011010110101000,
		32'b01110100000010110011011000000100,
		32'b01110011111000000011011001011111,
		32'b01110011101101010011011010111010,
		32'b01110011100010100011011100010100,
		32'b01110011010111110011011101101111,
		32'b01110011001100110011011111001010,
		32'b01110011000001110011100000100100,
		32'b01110010110110110011100001111110,
		32'b01110010101011110011100011011000,
		32'b01110010100000100011100100110010,
		32'b01110010010101010011100110001100,
		32'b01110010001001110011100111100110,
		32'b01110001111110100011101001000000,
		32'b01110001110011000011101010011001,
		32'b01110001100111100011101011110010,
		32'b01110001011011110011101101001100,
		32'b01110001010000010011101110100101,
		32'b01110001000100100011101111111101,
		32'b01110000111000100011110001010110,
		32'b01110000101100110011110010101111,
		32'b01110000100000110011110100000111,
		32'b01110000010100110011110101100000,
		32'b01110000001000110011110110111000,
		32'b01101111111100100011111000010000,
		32'b01101111110000010011111001101000,
		32'b01101111100100000011111010111111,
		32'b01101111010111110011111100010111,
		32'b01101111001011010011111101101110,
		32'b01101110111110110011111111000101,
		32'b01101110110010010100000000011101,
		32'b01101110100101100100000001110011,
		32'b01101110011000110100000011001010,
		32'b01101110001100000100000100100001,
		32'b01101101111111010100000101110111,
		32'b01101101110010100100000111001110,
		32'b01101101100101100100001000100100,
		32'b01101101011000100100001001111010,
		32'b01101101001011010100001011010000,
		32'b01101100111110010100001100100101,
		32'b01101100110001000100001101111011,
		32'b01101100100011110100001111010000,
		32'b01101100010110010100010000100101,
		32'b01101100001001000100010001111010,
		32'b01101011111011100100010011001111,
		32'b01101011101110000100010100100100,
		32'b01101011100000010100010101111000,
		32'b01101011010010100100010111001101,
		32'b01101011000100110100011000100001,
		32'b01101010110111000100011001110101,
		32'b01101010101001010100011011001001,
		32'b01101010011011010100011100011100,
		32'b01101010001101010100011101110000,
		32'b01101001111111010100011111000011,
		32'b01101001110001000100100000010110,
		32'b01101001100011000100100001101001,
		32'b01101001010100110100100010111100,
		32'b01101001000110010100100100001111,
		32'b01101000111000000100100101100001,
		32'b01101000101001100100100110110100,
		32'b01101000011011000100101000000110,
		32'b01101000001100100100101001011000,
		32'b01100111111101110100101010101001,
		32'b01100111101111010100101011111011,
		32'b01100111100000100100101101001100,
		32'b01100111010001100100101110011110,
		32'b01100111000010110100101111101111,
		32'b01100110110011110100110000111111,
		32'b01100110100100110100110010010000,
		32'b01100110010101110100110011100001,
		32'b01100110000110100100110100110001,
		32'b01100101110111010100110110000001,
		32'b01100101101000000100110111010001,
		32'b01100101011000110100111000100001,
		32'b01100101001001100100111001110000,
		32'b01100100111010000100111010111111,
		32'b01100100101010100100111100001111,
		32'b01100100011011000100111101011110,
		32'b01100100001011010100111110101100,
		32'b01100011111011110100111111111011,
		32'b01100011101100000101000001001001,
		32'b01100011011100010101000010010111,
		32'b01100011001100010101000011100101,
		32'b01100010111100100101000100110011,
		32'b01100010101100100101000110000001,
		32'b01100010011100010101000111001110,
		32'b01100010001100010101001000011100,
		32'b01100001111100010101001001101001,
		32'b01100001101100000101001010110101,
		32'b01100001011011110101001100000010,
		32'b01100001001011010101001101001110,
		32'b01100000111011000101001110011011,
		32'b01100000101010100101001111100111,
		32'b01100000011010000101010000110011,
		32'b01100000001001100101010001111110,
		32'b01011111111000110101010011001010,
		32'b01011111101000000101010100010101,
		32'b01011111010111100101010101100000,
		32'b01011111000110100101010110101011,
		32'b01011110110101110101010111110101,
		32'b01011110100100110101011001000000,
		32'b01011110010100000101011010001010,
		32'b01011110000010110101011011010100,
		32'b01011101110001110101011100011101,
		32'b01011101100000110101011101100111,
		32'b01011101001111100101011110110000,
		32'b01011100111110010101011111111001,
		32'b01011100101101000101100001000010,
		32'b01011100011011100101100010001011,
		32'b01011100001010010101100011010100,
		32'b01011011111000110101100100011100,
		32'b01011011100111010101100101100100,
		32'b01011011010101100101100110101100,
		32'b01011011000100000101100111110011,
		32'b01011010110010010101101000111011,
		32'b01011010100000100101101010000010,
		32'b01011010001110110101101011001001,
		32'b01011001111100110101101100010000,
		32'b01011001101011000101101101010110,
		32'b01011001011001000101101110011101,
		32'b01011001000111000101101111100011,
		32'b01011000110101000101110000101001,
		32'b01011000100010110101110001101110,
		32'b01011000010000100101110010110100,
		32'b01010111111110010101110011111001,
		32'b01010111101100000101110100111110,
		32'b01010111011001110101110110000011,
		32'b01010111000111010101110111000111,
		32'b01010110110101000101111000001011,
		32'b01010110100010100101111001010000,
		32'b01010110010000000101111010010011,
		32'b01010101111101010101111011010111,
		32'b01010101101010110101111100011010,
		32'b01010101011000000101111101011110,
		32'b01010101000101010101111110100000,
		32'b01010100110010100101111111100011,
		32'b01010100011111100110000000100110,
		32'b01010100001100110110000001101000,
		32'b01010011111001110110000010101010,
		32'b01010011100110110110000011101100,
		32'b01010011010011100110000100101101,
		32'b01010011000000100110000101101111,
		32'b01010010101101010110000110110000,
		32'b01010010011010010110000111110001,
		32'b01010010000111000110001000110001,
		32'b01010001110011100110001001110001,
		32'b01010001100000010110001010110010,
		32'b01010001001100110110001011110010,
		32'b01010000111001010110001100110001,
		32'b01010000100101110110001101110001,
		32'b01010000010010010110001110110000,
		32'b01001111111110110110001111101111,
		32'b01001111101011000110010000101101,
		32'b01001111010111100110010001101100,
		32'b01001111000011110110010010101010,
		32'b01001110101111110110010011101000,
		32'b01001110011100000110010100100110,
		32'b01001110001000010110010101100011,
		32'b01001101110100010110010110100000,
		32'b01001101100000010110010111011101,
		32'b01001101001100010110011000011010,
		32'b01001100111000010110011001010111,
		32'b01001100100100000110011010010011,
		32'b01001100001111110110011011001111,
		32'b01001011111011110110011100001011,
		32'b01001011100111100110011101000110,
		32'b01001011010011000110011110000010,
		32'b01001010111110110110011110111101,
		32'b01001010101010010110011111110111,
		32'b01001010010110000110100000110010,
		32'b01001010000001100110100001101100,
		32'b01001001101101000110100010100110,
		32'b01001001011000010110100011100000,
		32'b01001001000011110110100100011001,
		32'b01001000101111000110100101010011,
		32'b01001000011010010110100110001100,
		32'b01001000000101100110100111000100,
		32'b01000111110000110110100111111101,
		32'b01000111011100000110101000110101,
		32'b01000111000111000110101001101101,
		32'b01000110110010010110101010100101,
		32'b01000110011101010110101011011100,
		32'b01000110001000010110101100010011,
		32'b01000101110011010110101101001010,
		32'b01000101011110000110101110000001,
		32'b01000101001001000110101110111000,
		32'b01000100110011110110101111101110,
		32'b01000100011110100110110000100100,
		32'b01000100001001010110110001011001,
		32'b01000011110100000110110010001111,
		32'b01000011011110110110110011000100,
		32'b01000011001001010110110011111001,
		32'b01000010110100000110110100101101,
		32'b01000010011110100110110101100010,
		32'b01000010001001000110110110010110,
		32'b01000001110011100110110111001010,
		32'b01000001011101110110110111111101,
		32'b01000001001000010110111000110000,
		32'b01000000110010100110111001100011,
		32'b01000000011100110110111010010110,
		32'b01000000000111010110111011001001,
		32'b00111111110001010110111011111011,
		32'b00111111011011100110111100101101,
		32'b00111111000101110110111101011111,
		32'b00111110101111110110111110010000,
		32'b00111110011010000110111111000001,
		32'b00111110000100000110111111110010,
		32'b00111101101110000111000000100011,
		32'b00111101011000000111000001010011,
		32'b00111101000001110111000010000011,
		32'b00111100101011110111000010110011,
		32'b00111100010101100111000011100010,
		32'b00111011111111010111000100010010,
		32'b00111011101001010111000101000001,
		32'b00111011010011000111000101101111,
		32'b00111010111100100111000110011110,
		32'b00111010100110010111000111001100,
		32'b00111010010000000111000111111010,
		32'b00111001111001100111001000100111,
		32'b00111001100011000111001001010101,
		32'b00111001001100100111001010000010,
		32'b00111000110110000111001010101111,
		32'b00111000011111100111001011011011,
		32'b00111000001001000111001100000111,
		32'b00110111110010100111001100110011,
		32'b00110111011011110111001101011111,
		32'b00110111000101000111001110001010,
		32'b00110110101110100111001110110101,
		32'b00110110010111110111001111100000,
		32'b00110110000001000111010000001011,
		32'b00110101101010000111010000110101,
		32'b00110101010011010111010001011111,
		32'b00110100111100100111010010001001,
		32'b00110100100101100111010010110010,
		32'b00110100001110100111010011011011,
		32'b00110011110111100111010100000100,
		32'b00110011100000100111010100101101,
		32'b00110011001001100111010101010101,
		32'b00110010110010100111010101111101,
		32'b00110010011011100111010110100101,
		32'b00110010000100010111010111001100,
		32'b00110001101101010111010111110100,
		32'b00110001010110000111011000011011,
		32'b00110000111110110111011001000001,
		32'b00110000100111100111011001101000,
		32'b00110000010000010111011010001110,
		32'b00101111111001000111011010110011,
		32'b00101111100001110111011011011001,
		32'b00101111001010010111011011111110,
		32'b00101110110011000111011100100011,
		32'b00101110011011100111011101000111,
		32'b00101110000100010111011101101100,
		32'b00101101101100110111011110010000,
		32'b00101101010101010111011110110100,
		32'b00101100111101110111011111010111,
		32'b00101100100110000111011111111010,
		32'b00101100001110100111100000011101,
		32'b00101011110111000111100001000000,
		32'b00101011011111010111100001100010,
		32'b00101011000111110111100010000100,
		32'b00101010110000000111100010100110,
		32'b00101010011000010111100011000111,
		32'b00101010000000100111100011101000,
		32'b00101001101000110111100100001001,
		32'b00101001010001000111100100101010,
		32'b00101000111001010111100101001010,
		32'b00101000100001100111100101101010,
		32'b00101000001001100111100110001010,
		32'b00100111110001110111100110101001,
		32'b00100111011001110111100111001000,
		32'b00100111000001110111100111100111,
		32'b00100110101010000111101000000101,
		32'b00100110010010000111101000100100,
		32'b00100101111010000111101001000010,
		32'b00100101100010000111101001011111,
		32'b00100101001010000111101001111101,
		32'b00100100110001110111101010011010,
		32'b00100100011001110111101010110110,
		32'b00100100000001110111101011010011,
		32'b00100011101001100111101011101111,
		32'b00100011010001010111101100001011,
		32'b00100010111001010111101100100110,
		32'b00100010100001000111101101000010,
		32'b00100010001000110111101101011101,
		32'b00100001110000100111101101110111,
		32'b00100001011000010111101110010010,
		32'b00100001000000000111101110101100,
		32'b00100000100111110111101111000101,
		32'b00100000001111100111101111011111,
		32'b00011111110111000111101111111000,
		32'b00011111011110110111110000010001,
		32'b00011111000110010111110000101001,
		32'b00011110101110000111110001000010,
		32'b00011110010101100111110001011010,
		32'b00011101111101010111110001110001,
		32'b00011101100100110111110010001001,
		32'b00011101001100010111110010100000,
		32'b00011100110011110111110010110111,
		32'b00011100011011010111110011001101,
		32'b00011100000010110111110011100011,
		32'b00011011101010010111110011111001,
		32'b00011011010001110111110100001111,
		32'b00011010111001000111110100100100,
		32'b00011010100000100111110100111001,
		32'b00011010001000000111110101001110,
		32'b00011001101111010111110101100010,
		32'b00011001010110110111110101110110,
		32'b00011000111110000111110110001010,
		32'b00011000100101100111110110011101,
		32'b00011000001100110111110110110000,
		32'b00010111110100000111110111000011,
		32'b00010111011011010111110111010110,
		32'b00010111000010100111110111101000,
		32'b00010110101010000111110111111010,
		32'b00010110010001010111111000001100,
		32'b00010101111000100111111000011101,
		32'b00010101011111110111111000101110,
		32'b00010101000110110111111000111111,
		32'b00010100101110000111111001001111,
		32'b00010100010101010111111001011111,
		32'b00010011111100100111111001101111,
		32'b00010011100011100111111001111111,
		32'b00010011001010110111111010001110,
		32'b00010010110010000111111010011101,
		32'b00010010011001000111111010101011,
		32'b00010010000000010111111010111010,
		32'b00010001100111010111111011001000,
		32'b00010001001110010111111011010101,
		32'b00010000110101100111111011100011,
		32'b00010000011100100111111011110000,
		32'b00010000000011100111111011111101,
		32'b00001111101010110111111100001001,
		32'b00001111010001110111111100010101,
		32'b00001110111000110111111100100001,
		32'b00001110011111110111111100101101,
		32'b00001110000110110111111100111000,
		32'b00001101101101110111111101000011,
		32'b00001101010100110111111101001101,
		32'b00001100111011110111111101011000,
		32'b00001100100010110111111101100010,
		32'b00001100001001110111111101101011,
		32'b00001011110000110111111101110101,
		32'b00001011010111110111111101111110,
		32'b00001010111110110111111110000111,
		32'b00001010100101110111111110001111,
		32'b00001010001100110111111110010111,
		32'b00001001110011100111111110011111,
		32'b00001001011010100111111110100111,
		32'b00001001000001100111111110101110,
		32'b00001000101000100111111110110101,
		32'b00001000001111010111111110111100,
		32'b00000111110110010111111111000010,
		32'b00000111011101010111111111001000,
		32'b00000111000100000111111111001110,
		32'b00000110101011000111111111010011,
		32'b00000110010001110111111111011000,
		32'b00000101111000110111111111011101,
		32'b00000101011111110111111111100001,
		32'b00000101000110100111111111100101,
		32'b00000100101101100111111111101001,
		32'b00000100010100010111111111101101,
		32'b00000011111011010111111111110000,
		32'b00000011100010000111111111110011,
		32'b00000011001001000111111111110110,
		32'b00000010101111110111111111111000,
		32'b00000010010110110111111111111010,
		32'b00000001111101100111111111111100,
		32'b00000001100100100111111111111101,
		32'b00000001001011010111111111111110,
		32'b00000000110010010111111111111111,
		32'b00000000011001000111111111111111,
		32'b00000000000000000111111111111111,
		32'b10000000011001000111111111111111,
		32'b10000000110010010111111111111111,
		32'b10000001001011010111111111111110,
		32'b10000001100100100111111111111101,
		32'b10000001111101100111111111111100,
		32'b10000010010110110111111111111010,
		32'b10000010101111110111111111111000,
		32'b10000011001001000111111111110110,
		32'b10000011100010000111111111110011,
		32'b10000011111011010111111111110000,
		32'b10000100010100010111111111101101,
		32'b10000100101101100111111111101001,
		32'b10000101000110100111111111100101,
		32'b10000101011111110111111111100001,
		32'b10000101111000110111111111011101,
		32'b10000110010001110111111111011000,
		32'b10000110101011000111111111010011,
		32'b10000111000100000111111111001110,
		32'b10000111011101010111111111001000,
		32'b10000111110110010111111111000010,
		32'b10001000001111010111111110111100,
		32'b10001000101000100111111110110101,
		32'b10001001000001100111111110101110,
		32'b10001001011010100111111110100111,
		32'b10001001110011100111111110011111,
		32'b10001010001100110111111110010111,
		32'b10001010100101110111111110001111,
		32'b10001010111110110111111110000111,
		32'b10001011010111110111111101111110,
		32'b10001011110000110111111101110101,
		32'b10001100001001110111111101101011,
		32'b10001100100010110111111101100010,
		32'b10001100111011110111111101011000,
		32'b10001101010100110111111101001101,
		32'b10001101101101110111111101000011,
		32'b10001110000110110111111100111000,
		32'b10001110011111110111111100101101,
		32'b10001110111000110111111100100001,
		32'b10001111010001110111111100010101,
		32'b10001111101010110111111100001001,
		32'b10010000000011100111111011111101,
		32'b10010000011100100111111011110000,
		32'b10010000110101100111111011100011,
		32'b10010001001110010111111011010101,
		32'b10010001100111010111111011001000,
		32'b10010010000000010111111010111010,
		32'b10010010011001000111111010101011,
		32'b10010010110010000111111010011101,
		32'b10010011001010110111111010001110,
		32'b10010011100011100111111001111111,
		32'b10010011111100100111111001101111,
		32'b10010100010101010111111001011111,
		32'b10010100101110000111111001001111,
		32'b10010101000110110111111000111111,
		32'b10010101011111110111111000101110,
		32'b10010101111000100111111000011101,
		32'b10010110010001010111111000001100,
		32'b10010110101010000111110111111010,
		32'b10010111000010100111110111101000,
		32'b10010111011011010111110111010110,
		32'b10010111110100000111110111000011,
		32'b10011000001100110111110110110000,
		32'b10011000100101100111110110011101,
		32'b10011000111110000111110110001010,
		32'b10011001010110110111110101110110,
		32'b10011001101111010111110101100010,
		32'b10011010001000000111110101001110,
		32'b10011010100000100111110100111001,
		32'b10011010111001000111110100100100,
		32'b10011011010001110111110100001111,
		32'b10011011101010010111110011111001,
		32'b10011100000010110111110011100011,
		32'b10011100011011010111110011001101,
		32'b10011100110011110111110010110111,
		32'b10011101001100010111110010100000,
		32'b10011101100100110111110010001001,
		32'b10011101111101010111110001110001,
		32'b10011110010101100111110001011010,
		32'b10011110101110000111110001000010,
		32'b10011111000110010111110000101001,
		32'b10011111011110110111110000010001,
		32'b10011111110111000111101111111000,
		32'b10100000001111100111101111011111,
		32'b10100000100111110111101111000101,
		32'b10100001000000000111101110101100,
		32'b10100001011000010111101110010010,
		32'b10100001110000100111101101110111,
		32'b10100010001000110111101101011101,
		32'b10100010100001000111101101000010,
		32'b10100010111001010111101100100110,
		32'b10100011010001010111101100001011,
		32'b10100011101001100111101011101111,
		32'b10100100000001110111101011010011,
		32'b10100100011001110111101010110110,
		32'b10100100110001110111101010011010,
		32'b10100101001010000111101001111101,
		32'b10100101100010000111101001011111,
		32'b10100101111010000111101001000010,
		32'b10100110010010000111101000100100,
		32'b10100110101010000111101000000101,
		32'b10100111000001110111100111100111,
		32'b10100111011001110111100111001000,
		32'b10100111110001110111100110101001,
		32'b10101000001001100111100110001010,
		32'b10101000100001100111100101101010,
		32'b10101000111001010111100101001010,
		32'b10101001010001000111100100101010,
		32'b10101001101000110111100100001001,
		32'b10101010000000100111100011101000,
		32'b10101010011000010111100011000111,
		32'b10101010110000000111100010100110,
		32'b10101011000111110111100010000100,
		32'b10101011011111010111100001100010,
		32'b10101011110111000111100001000000,
		32'b10101100001110100111100000011101,
		32'b10101100100110000111011111111010,
		32'b10101100111101110111011111010111,
		32'b10101101010101010111011110110100,
		32'b10101101101100110111011110010000,
		32'b10101110000100010111011101101100,
		32'b10101110011011100111011101000111,
		32'b10101110110011000111011100100011,
		32'b10101111001010010111011011111110,
		32'b10101111100001110111011011011001,
		32'b10101111111001000111011010110011,
		32'b10110000010000010111011010001110,
		32'b10110000100111100111011001101000,
		32'b10110000111110110111011001000001,
		32'b10110001010110000111011000011011,
		32'b10110001101101010111010111110100,
		32'b10110010000100010111010111001100,
		32'b10110010011011100111010110100101,
		32'b10110010110010100111010101111101,
		32'b10110011001001100111010101010101,
		32'b10110011100000100111010100101101,
		32'b10110011110111100111010100000100,
		32'b10110100001110100111010011011011,
		32'b10110100100101100111010010110010,
		32'b10110100111100100111010010001001,
		32'b10110101010011010111010001011111,
		32'b10110101101010000111010000110101,
		32'b10110110000001000111010000001011,
		32'b10110110010111110111001111100000,
		32'b10110110101110100111001110110101,
		32'b10110111000101000111001110001010,
		32'b10110111011011110111001101011111,
		32'b10110111110010100111001100110011,
		32'b10111000001001000111001100000111,
		32'b10111000011111100111001011011011,
		32'b10111000110110000111001010101111,
		32'b10111001001100100111001010000010,
		32'b10111001100011000111001001010101,
		32'b10111001111001100111001000100111,
		32'b10111010010000000111000111111010,
		32'b10111010100110010111000111001100,
		32'b10111010111100100111000110011110,
		32'b10111011010011000111000101101111,
		32'b10111011101001010111000101000001,
		32'b10111011111111010111000100010010,
		32'b10111100010101100111000011100010,
		32'b10111100101011110111000010110011,
		32'b10111101000001110111000010000011,
		32'b10111101011000000111000001010011,
		32'b10111101101110000111000000100011,
		32'b10111110000100000110111111110010,
		32'b10111110011010000110111111000001,
		32'b10111110101111110110111110010000,
		32'b10111111000101110110111101011111,
		32'b10111111011011100110111100101101,
		32'b10111111110001010110111011111011,
		32'b11000000000111010110111011001001,
		32'b11000000011100110110111010010110,
		32'b11000000110010100110111001100011,
		32'b11000001001000010110111000110000,
		32'b11000001011101110110110111111101,
		32'b11000001110011100110110111001010,
		32'b11000010001001000110110110010110,
		32'b11000010011110100110110101100010,
		32'b11000010110100000110110100101101,
		32'b11000011001001010110110011111001,
		32'b11000011011110110110110011000100,
		32'b11000011110100000110110010001111,
		32'b11000100001001010110110001011001,
		32'b11000100011110100110110000100100,
		32'b11000100110011110110101111101110,
		32'b11000101001001000110101110111000,
		32'b11000101011110000110101110000001,
		32'b11000101110011010110101101001010,
		32'b11000110001000010110101100010011,
		32'b11000110011101010110101011011100,
		32'b11000110110010010110101010100101,
		32'b11000111000111000110101001101101,
		32'b11000111011100000110101000110101,
		32'b11000111110000110110100111111101,
		32'b11001000000101100110100111000100,
		32'b11001000011010010110100110001100,
		32'b11001000101111000110100101010011,
		32'b11001001000011110110100100011001,
		32'b11001001011000010110100011100000,
		32'b11001001101101000110100010100110,
		32'b11001010000001100110100001101100,
		32'b11001010010110000110100000110010,
		32'b11001010101010010110011111110111,
		32'b11001010111110110110011110111101,
		32'b11001011010011000110011110000010,
		32'b11001011100111100110011101000110,
		32'b11001011111011110110011100001011,
		32'b11001100001111110110011011001111,
		32'b11001100100100000110011010010011,
		32'b11001100111000010110011001010111,
		32'b11001101001100010110011000011010,
		32'b11001101100000010110010111011101,
		32'b11001101110100010110010110100000,
		32'b11001110001000010110010101100011,
		32'b11001110011100000110010100100110,
		32'b11001110101111110110010011101000,
		32'b11001111000011110110010010101010,
		32'b11001111010111100110010001101100,
		32'b11001111101011000110010000101101,
		32'b11001111111110110110001111101111,
		32'b11010000010010010110001110110000,
		32'b11010000100101110110001101110001,
		32'b11010000111001010110001100110001,
		32'b11010001001100110110001011110010,
		32'b11010001100000010110001010110010,
		32'b11010001110011100110001001110001,
		32'b11010010000111000110001000110001,
		32'b11010010011010010110000111110001,
		32'b11010010101101010110000110110000,
		32'b11010011000000100110000101101111,
		32'b11010011010011100110000100101101,
		32'b11010011100110110110000011101100,
		32'b11010011111001110110000010101010,
		32'b11010100001100110110000001101000,
		32'b11010100011111100110000000100110,
		32'b11010100110010100101111111100011,
		32'b11010101000101010101111110100000,
		32'b11010101011000000101111101011110,
		32'b11010101101010110101111100011010,
		32'b11010101111101010101111011010111,
		32'b11010110010000000101111010010011,
		32'b11010110100010100101111001010000,
		32'b11010110110101000101111000001011,
		32'b11010111000111010101110111000111,
		32'b11010111011001110101110110000011,
		32'b11010111101100000101110100111110,
		32'b11010111111110010101110011111001,
		32'b11011000010000100101110010110100,
		32'b11011000100010110101110001101110,
		32'b11011000110101000101110000101001,
		32'b11011001000111000101101111100011,
		32'b11011001011001000101101110011101,
		32'b11011001101011000101101101010110,
		32'b11011001111100110101101100010000,
		32'b11011010001110110101101011001001,
		32'b11011010100000100101101010000010,
		32'b11011010110010010101101000111011,
		32'b11011011000100000101100111110011,
		32'b11011011010101100101100110101100,
		32'b11011011100111010101100101100100,
		32'b11011011111000110101100100011100,
		32'b11011100001010010101100011010100,
		32'b11011100011011100101100010001011,
		32'b11011100101101000101100001000010,
		32'b11011100111110010101011111111001,
		32'b11011101001111100101011110110000,
		32'b11011101100000110101011101100111,
		32'b11011101110001110101011100011101,
		32'b11011110000010110101011011010100,
		32'b11011110010100000101011010001010,
		32'b11011110100100110101011001000000,
		32'b11011110110101110101010111110101,
		32'b11011111000110100101010110101011,
		32'b11011111010111100101010101100000,
		32'b11011111101000000101010100010101,
		32'b11011111111000110101010011001010,
		32'b11100000001001100101010001111110,
		32'b11100000011010000101010000110011,
		32'b11100000101010100101001111100111,
		32'b11100000111011000101001110011011,
		32'b11100001001011010101001101001110,
		32'b11100001011011110101001100000010,
		32'b11100001101100000101001010110101,
		32'b11100001111100010101001001101001,
		32'b11100010001100010101001000011100,
		32'b11100010011100010101000111001110,
		32'b11100010101100100101000110000001,
		32'b11100010111100100101000100110011,
		32'b11100011001100010101000011100101,
		32'b11100011011100010101000010010111,
		32'b11100011101100000101000001001001,
		32'b11100011111011110100111111111011,
		32'b11100100001011010100111110101100,
		32'b11100100011011000100111101011110,
		32'b11100100101010100100111100001111,
		32'b11100100111010000100111010111111,
		32'b11100101001001100100111001110000,
		32'b11100101011000110100111000100001,
		32'b11100101101000000100110111010001,
		32'b11100101110111010100110110000001,
		32'b11100110000110100100110100110001,
		32'b11100110010101110100110011100001,
		32'b11100110100100110100110010010000,
		32'b11100110110011110100110000111111,
		32'b11100111000010110100101111101111,
		32'b11100111010001100100101110011110,
		32'b11100111100000100100101101001100,
		32'b11100111101111010100101011111011,
		32'b11100111111101110100101010101001,
		32'b11101000001100100100101001011000,
		32'b11101000011011000100101000000110,
		32'b11101000101001100100100110110100,
		32'b11101000111000000100100101100001,
		32'b11101001000110010100100100001111,
		32'b11101001010100110100100010111100,
		32'b11101001100011000100100001101001,
		32'b11101001110001000100100000010110,
		32'b11101001111111010100011111000011,
		32'b11101010001101010100011101110000,
		32'b11101010011011010100011100011100,
		32'b11101010101001010100011011001001,
		32'b11101010110111000100011001110101,
		32'b11101011000100110100011000100001,
		32'b11101011010010100100010111001101,
		32'b11101011100000010100010101111000,
		32'b11101011101110000100010100100100,
		32'b11101011111011100100010011001111,
		32'b11101100001001000100010001111010,
		32'b11101100010110010100010000100101,
		32'b11101100100011110100001111010000,
		32'b11101100110001000100001101111011,
		32'b11101100111110010100001100100101,
		32'b11101101001011010100001011010000,
		32'b11101101011000100100001001111010,
		32'b11101101100101100100001000100100,
		32'b11101101110010100100000111001110,
		32'b11101101111111010100000101110111,
		32'b11101110001100000100000100100001,
		32'b11101110011000110100000011001010,
		32'b11101110100101100100000001110011,
		32'b11101110110010010100000000011101,
		32'b11101110111110110011111111000101,
		32'b11101111001011010011111101101110,
		32'b11101111010111110011111100010111,
		32'b11101111100100000011111010111111,
		32'b11101111110000010011111001101000,
		32'b11101111111100100011111000010000,
		32'b11110000001000110011110110111000,
		32'b11110000010100110011110101100000,
		32'b11110000100000110011110100000111,
		32'b11110000101100110011110010101111,
		32'b11110000111000100011110001010110,
		32'b11110001000100100011101111111101,
		32'b11110001010000010011101110100101,
		32'b11110001011011110011101101001100,
		32'b11110001100111100011101011110010,
		32'b11110001110011000011101010011001,
		32'b11110001111110100011101001000000,
		32'b11110010001001110011100111100110,
		32'b11110010010101010011100110001100,
		32'b11110010100000100011100100110010,
		32'b11110010101011110011100011011000,
		32'b11110010110110110011100001111110,
		32'b11110011000001110011100000100100,
		32'b11110011001100110011011111001010,
		32'b11110011010111110011011101101111,
		32'b11110011100010100011011100010100,
		32'b11110011101101010011011010111010,
		32'b11110011111000000011011001011111,
		32'b11110100000010110011011000000100,
		32'b11110100001101010011010110101000,
		32'b11110100010111110011010101001101,
		32'b11110100100010010011010011110010,
		32'b11110100101100100011010010010110,
		32'b11110100110110110011010000111010,
		32'b11110101000001000011001111011110,
		32'b11110101001011010011001110000010,
		32'b11110101010101010011001100100110,
		32'b11110101011111010011001011001010,
		32'b11110101101001010011001001101110,
		32'b11110101110011000011001000010001,
		32'b11110101111101000011000110110101,
		32'b11110110000110110011000101011000,
		32'b11110110010000010011000011111011,
		32'b11110110011010000011000010011110,
		32'b11110110100011100011000001000001,
		32'b11110110101100110010111111100100,
		32'b11110110110110010010111110000111,
		32'b11110110111111100010111100101001,
		32'b11110111001000110010111011001100,
		32'b11110111010001110010111001101110,
		32'b11110111011011000010111000010001,
		32'b11110111100100000010110110110011,
		32'b11110111101101000010110101010101,
		32'b11110111110101110010110011110111,
		32'b11110111111110100010110010011000,
		32'b11111000000111010010110000111010,
		32'b11111000010000000010101111011100,
		32'b11111000011000100010101101111101,
		32'b11111000100001000010101100011111,
		32'b11111000101001100010101011000000,
		32'b11111000110001110010101001100001,
		32'b11111000111010000010101000000010,
		32'b11111001000010010010100110100011,
		32'b11111001001010100010100101000100,
		32'b11111001010010100010100011100101,
		32'b11111001011010100010100010000110,
		32'b11111001100010100010100000100110,
		32'b11111001101010010010011111000111,
		32'b11111001110010000010011101100111,
		32'b11111001111001110010011100000111,
		32'b11111010000001010010011010101000,
		32'b11111010001001000010011001001000,
		32'b11111010010000100010010111101000,
		32'b11111010010111110010010110001000,
		32'b11111010011111010010010100101000,
		32'b11111010100110100010010011000111,
		32'b11111010101101100010010001100111,
		32'b11111010110100110010010000000111,
		32'b11111010111011110010001110100110,
		32'b11111011000010110010001101000101,
		32'b11111011001001100010001011100101,
		32'b11111011010000100010001010000100,
		32'b11111011010111010010001000100011,
		32'b11111011011101110010000111000010,
		32'b11111011100100100010000101100001,
		32'b11111011101011000010000100000000,
		32'b11111011110001010010000010011111,
		32'b11111011110111110010000000111110,
		32'b11111011111110000001111111011100,
		32'b11111100000100010001111101111011,
		32'b11111100001010010001111100011001,
		32'b11111100010000100001111010111000,
		32'b11111100010110100001111001010110,
		32'b11111100011100010001110111110101,
		32'b11111100100010010001110110010011,
		32'b11111100101000000001110100110001,
		32'b11111100101101110001110011001111,
		32'b11111100110011010001110001101101,
		32'b11111100111000110001110000001011,
		32'b11111100111110010001101110101001,
		32'b11111101000011110001101101000111,
		32'b11111101001001000001101011100100,
		32'b11111101001110010001101010000010,
		32'b11111101010011100001101000100000,
		32'b11111101011000100001100110111101,
		32'b11111101011101100001100101011011,
		32'b11111101100010100001100011111000,
		32'b11111101100111010001100010010110,
		32'b11111101101100000001100000110011,
		32'b11111101110000110001011111010000,
		32'b11111101110101100001011101101101,
		32'b11111101111010000001011100001010,
		32'b11111101111110100001011010101000,
		32'b11111110000011000001011001000101,
		32'b11111110000111010001010111100010,
		32'b11111110001011100001010101111111,
		32'b11111110001111110001010100011011,
		32'b11111110010011110001010010111000,
		32'b11111110010111110001010001010101,
		32'b11111110011011110001001111110010,
		32'b11111110011111110001001110001110,
		32'b11111110100011100001001100101011,
		32'b11111110100111010001001011001000,
		32'b11111110101010110001001001100100,
		32'b11111110101110100001001000000001,
		32'b11111110110010000001000110011101,
		32'b11111110110101010001000100111001,
		32'b11111110111000110001000011010110,
		32'b11111110111100000001000001110010,
		32'b11111110111111010001000000001110,
		32'b11111111000010010000111110101011,
		32'b11111111000101010000111101000111,
		32'b11111111001000010000111011100011,
		32'b11111111001011010000111001111111,
		32'b11111111001110000000111000011011,
		32'b11111111010000110000110110110111,
		32'b11111111010011010000110101010011,
		32'b11111111010110000000110011101111,
		32'b11111111011000100000110010001011,
		32'b11111111011010110000110000100111,
		32'b11111111011101010000101111000011,
		32'b11111111011111100000101101011111,
		32'b11111111100001110000101011111011,
		32'b11111111100011110000101010010111,
		32'b11111111100101110000101000110011,
		32'b11111111100111110000100111001110,
		32'b11111111101001110000100101101010,
		32'b11111111101011100000100100000110,
		32'b11111111101101010000100010100010,
		32'b11111111101111000000100000111101,
		32'b11111111110000100000011111011001,
		32'b11111111110010000000011101110101,
		32'b11111111110011100000011100010000,
		32'b11111111110100110000011010101100,
		32'b11111111110110000000011001000111,
		32'b11111111110111010000010111100011,
		32'b11111111111000010000010101111111,
		32'b11111111111001010000010100011010,
		32'b11111111111010010000010010110110,
		32'b11111111111011010000010001010001,
		32'b11111111111100000000001111101101,
		32'b11111111111100110000001110001000,
		32'b11111111111101100000001100100100,
		32'b11111111111110000000001010111111,
		32'b11111111111110100000001001011011,
		32'b11111111111111000000000111110110,
		32'b11111111111111010000000110010010,
		32'b11111111111111100000000100101101,
		32'b11111111111111110000000011001001,
		32'b11111111111111110000000001100100,
		32'b11111111111111110000000000000000,
		32'b11111111111111111000000001100100,
		32'b11111111111111111000000011001001,
		32'b11111111111111101000000100101101,
		32'b11111111111111011000000110010010,
		32'b11111111111111001000000111110110,
		32'b11111111111110101000001001011011,
		32'b11111111111110001000001010111111,
		32'b11111111111101101000001100100100,
		32'b11111111111100111000001110001000,
		32'b11111111111100001000001111101101,
		32'b11111111111011011000010001010001,
		32'b11111111111010011000010010110110,
		32'b11111111111001011000010100011010,
		32'b11111111111000011000010101111111,
		32'b11111111110111011000010111100011,
		32'b11111111110110001000011001000111,
		32'b11111111110100111000011010101100,
		32'b11111111110011101000011100010000,
		32'b11111111110010001000011101110101,
		32'b11111111110000101000011111011001,
		32'b11111111101111001000100000111101,
		32'b11111111101101011000100010100010,
		32'b11111111101011101000100100000110,
		32'b11111111101001111000100101101010,
		32'b11111111100111111000100111001110,
		32'b11111111100101111000101000110011,
		32'b11111111100011111000101010010111,
		32'b11111111100001111000101011111011,
		32'b11111111011111101000101101011111,
		32'b11111111011101011000101111000011,
		32'b11111111011010111000110000100111,
		32'b11111111011000101000110010001011,
		32'b11111111010110001000110011101111,
		32'b11111111010011011000110101010011,
		32'b11111111010000111000110110110111,
		32'b11111111001110001000111000011011,
		32'b11111111001011011000111001111111,
		32'b11111111001000011000111011100011,
		32'b11111111000101011000111101000111,
		32'b11111111000010011000111110101011,
		32'b11111110111111011001000000001110,
		32'b11111110111100001001000001110010,
		32'b11111110111000111001000011010110,
		32'b11111110110101011001000100111001,
		32'b11111110110010001001000110011101,
		32'b11111110101110101001001000000001,
		32'b11111110101010111001001001100100,
		32'b11111110100111011001001011001000,
		32'b11111110100011101001001100101011,
		32'b11111110011111111001001110001110,
		32'b11111110011011111001001111110010,
		32'b11111110010111111001010001010101,
		32'b11111110010011111001010010111000,
		32'b11111110001111111001010100011011,
		32'b11111110001011101001010101111111,
		32'b11111110000111011001010111100010,
		32'b11111110000011001001011001000101,
		32'b11111101111110101001011010101000,
		32'b11111101111010001001011100001010,
		32'b11111101110101101001011101101101,
		32'b11111101110000111001011111010000,
		32'b11111101101100001001100000110011,
		32'b11111101100111011001100010010110,
		32'b11111101100010101001100011111000,
		32'b11111101011101101001100101011011,
		32'b11111101011000101001100110111101,
		32'b11111101010011101001101000100000,
		32'b11111101001110011001101010000010,
		32'b11111101001001001001101011100100,
		32'b11111101000011111001101101000111,
		32'b11111100111110011001101110101001,
		32'b11111100111000111001110000001011,
		32'b11111100110011011001110001101101,
		32'b11111100101101111001110011001111,
		32'b11111100101000001001110100110001,
		32'b11111100100010011001110110010011,
		32'b11111100011100011001110111110101,
		32'b11111100010110101001111001010110,
		32'b11111100010000101001111010111000,
		32'b11111100001010011001111100011001,
		32'b11111100000100011001111101111011,
		32'b11111011111110001001111111011100,
		32'b11111011110111111010000000111110,
		32'b11111011110001011010000010011111,
		32'b11111011101011001010000100000000,
		32'b11111011100100101010000101100001,
		32'b11111011011101111010000111000010,
		32'b11111011010111011010001000100011,
		32'b11111011010000101010001010000100,
		32'b11111011001001101010001011100101,
		32'b11111011000010111010001101000101,
		32'b11111010111011111010001110100110,
		32'b11111010110100111010010000000111,
		32'b11111010101101101010010001100111,
		32'b11111010100110101010010011000111,
		32'b11111010011111011010010100101000,
		32'b11111010010111111010010110001000,
		32'b11111010010000101010010111101000,
		32'b11111010001001001010011001001000,
		32'b11111010000001011010011010101000,
		32'b11111001111001111010011100000111,
		32'b11111001110010001010011101100111,
		32'b11111001101010011010011111000111,
		32'b11111001100010101010100000100110,
		32'b11111001011010101010100010000110,
		32'b11111001010010101010100011100101,
		32'b11111001001010101010100101000100,
		32'b11111001000010011010100110100011,
		32'b11111000111010001010101000000010,
		32'b11111000110001111010101001100001,
		32'b11111000101001101010101011000000,
		32'b11111000100001001010101100011111,
		32'b11111000011000101010101101111101,
		32'b11111000010000001010101111011100,
		32'b11111000000111011010110000111010,
		32'b11110111111110101010110010011000,
		32'b11110111110101111010110011110111,
		32'b11110111101101001010110101010101,
		32'b11110111100100001010110110110011,
		32'b11110111011011001010111000010001,
		32'b11110111010001111010111001101110,
		32'b11110111001000111010111011001100,
		32'b11110110111111101010111100101001,
		32'b11110110110110011010111110000111,
		32'b11110110101100111010111111100100,
		32'b11110110100011101011000001000001,
		32'b11110110011010001011000010011110,
		32'b11110110010000011011000011111011,
		32'b11110110000110111011000101011000,
		32'b11110101111101001011000110110101,
		32'b11110101110011001011001000010001,
		32'b11110101101001011011001001101110,
		32'b11110101011111011011001011001010,
		32'b11110101010101011011001100100110,
		32'b11110101001011011011001110000010,
		32'b11110101000001001011001111011110,
		32'b11110100110110111011010000111010,
		32'b11110100101100101011010010010110,
		32'b11110100100010011011010011110010,
		32'b11110100010111111011010101001101,
		32'b11110100001101011011010110101000,
		32'b11110100000010111011011000000100,
		32'b11110011111000001011011001011111,
		32'b11110011101101011011011010111010,
		32'b11110011100010101011011100010100,
		32'b11110011010111111011011101101111,
		32'b11110011001100111011011111001010,
		32'b11110011000001111011100000100100,
		32'b11110010110110111011100001111110,
		32'b11110010101011111011100011011000,
		32'b11110010100000101011100100110010,
		32'b11110010010101011011100110001100,
		32'b11110010001001111011100111100110,
		32'b11110001111110101011101001000000,
		32'b11110001110011001011101010011001,
		32'b11110001100111101011101011110010,
		32'b11110001011011111011101101001100,
		32'b11110001010000011011101110100101,
		32'b11110001000100101011101111111101,
		32'b11110000111000101011110001010110,
		32'b11110000101100111011110010101111,
		32'b11110000100000111011110100000111,
		32'b11110000010100111011110101100000,
		32'b11110000001000111011110110111000,
		32'b11101111111100101011111000010000,
		32'b11101111110000011011111001101000,
		32'b11101111100100001011111010111111,
		32'b11101111010111111011111100010111,
		32'b11101111001011011011111101101110,
		32'b11101110111110111011111111000101,
		32'b11101110110010011100000000011101,
		32'b11101110100101101100000001110011,
		32'b11101110011000111100000011001010,
		32'b11101110001100001100000100100001,
		32'b11101101111111011100000101110111,
		32'b11101101110010101100000111001110,
		32'b11101101100101101100001000100100,
		32'b11101101011000101100001001111010,
		32'b11101101001011011100001011010000,
		32'b11101100111110011100001100100101,
		32'b11101100110001001100001101111011,
		32'b11101100100011111100001111010000,
		32'b11101100010110011100010000100101,
		32'b11101100001001001100010001111010,
		32'b11101011111011101100010011001111,
		32'b11101011101110001100010100100100,
		32'b11101011100000011100010101111000,
		32'b11101011010010101100010111001101,
		32'b11101011000100111100011000100001,
		32'b11101010110111001100011001110101,
		32'b11101010101001011100011011001001,
		32'b11101010011011011100011100011100,
		32'b11101010001101011100011101110000,
		32'b11101001111111011100011111000011,
		32'b11101001110001001100100000010110,
		32'b11101001100011001100100001101001,
		32'b11101001010100111100100010111100,
		32'b11101001000110011100100100001111,
		32'b11101000111000001100100101100001,
		32'b11101000101001101100100110110100,
		32'b11101000011011001100101000000110,
		32'b11101000001100101100101001011000,
		32'b11100111111101111100101010101001,
		32'b11100111101111011100101011111011,
		32'b11100111100000101100101101001100,
		32'b11100111010001101100101110011110,
		32'b11100111000010111100101111101111,
		32'b11100110110011111100110000111111,
		32'b11100110100100111100110010010000,
		32'b11100110010101111100110011100001,
		32'b11100110000110101100110100110001,
		32'b11100101110111011100110110000001,
		32'b11100101101000001100110111010001,
		32'b11100101011000111100111000100001,
		32'b11100101001001101100111001110000,
		32'b11100100111010001100111010111111,
		32'b11100100101010101100111100001111,
		32'b11100100011011001100111101011110,
		32'b11100100001011011100111110101100,
		32'b11100011111011111100111111111011,
		32'b11100011101100001101000001001001,
		32'b11100011011100011101000010010111,
		32'b11100011001100011101000011100101,
		32'b11100010111100101101000100110011,
		32'b11100010101100101101000110000001,
		32'b11100010011100011101000111001110,
		32'b11100010001100011101001000011100,
		32'b11100001111100011101001001101001,
		32'b11100001101100001101001010110101,
		32'b11100001011011111101001100000010,
		32'b11100001001011011101001101001110,
		32'b11100000111011001101001110011011,
		32'b11100000101010101101001111100111,
		32'b11100000011010001101010000110011,
		32'b11100000001001101101010001111110,
		32'b11011111111000111101010011001010,
		32'b11011111101000001101010100010101,
		32'b11011111010111101101010101100000,
		32'b11011111000110101101010110101011,
		32'b11011110110101111101010111110101,
		32'b11011110100100111101011001000000,
		32'b11011110010100001101011010001010,
		32'b11011110000010111101011011010100,
		32'b11011101110001111101011100011101,
		32'b11011101100000111101011101100111,
		32'b11011101001111101101011110110000,
		32'b11011100111110011101011111111001,
		32'b11011100101101001101100001000010,
		32'b11011100011011101101100010001011,
		32'b11011100001010011101100011010100,
		32'b11011011111000111101100100011100,
		32'b11011011100111011101100101100100,
		32'b11011011010101101101100110101100,
		32'b11011011000100001101100111110011,
		32'b11011010110010011101101000111011,
		32'b11011010100000101101101010000010,
		32'b11011010001110111101101011001001,
		32'b11011001111100111101101100010000,
		32'b11011001101011001101101101010110,
		32'b11011001011001001101101110011101,
		32'b11011001000111001101101111100011,
		32'b11011000110101001101110000101001,
		32'b11011000100010111101110001101110,
		32'b11011000010000101101110010110100,
		32'b11010111111110011101110011111001,
		32'b11010111101100001101110100111110,
		32'b11010111011001111101110110000011,
		32'b11010111000111011101110111000111,
		32'b11010110110101001101111000001011,
		32'b11010110100010101101111001010000,
		32'b11010110010000001101111010010011,
		32'b11010101111101011101111011010111,
		32'b11010101101010111101111100011010,
		32'b11010101011000001101111101011110,
		32'b11010101000101011101111110100000,
		32'b11010100110010101101111111100011,
		32'b11010100011111101110000000100110,
		32'b11010100001100111110000001101000,
		32'b11010011111001111110000010101010,
		32'b11010011100110111110000011101100,
		32'b11010011010011101110000100101101,
		32'b11010011000000101110000101101111,
		32'b11010010101101011110000110110000,
		32'b11010010011010011110000111110001,
		32'b11010010000111001110001000110001,
		32'b11010001110011101110001001110001,
		32'b11010001100000011110001010110010,
		32'b11010001001100111110001011110010,
		32'b11010000111001011110001100110001,
		32'b11010000100101111110001101110001,
		32'b11010000010010011110001110110000,
		32'b11001111111110111110001111101111,
		32'b11001111101011001110010000101101,
		32'b11001111010111101110010001101100,
		32'b11001111000011111110010010101010,
		32'b11001110101111111110010011101000,
		32'b11001110011100001110010100100110,
		32'b11001110001000011110010101100011,
		32'b11001101110100011110010110100000,
		32'b11001101100000011110010111011101,
		32'b11001101001100011110011000011010,
		32'b11001100111000011110011001010111,
		32'b11001100100100001110011010010011,
		32'b11001100001111111110011011001111,
		32'b11001011111011111110011100001011,
		32'b11001011100111101110011101000110,
		32'b11001011010011001110011110000010,
		32'b11001010111110111110011110111101,
		32'b11001010101010011110011111110111,
		32'b11001010010110001110100000110010,
		32'b11001010000001101110100001101100,
		32'b11001001101101001110100010100110,
		32'b11001001011000011110100011100000,
		32'b11001001000011111110100100011001,
		32'b11001000101111001110100101010011,
		32'b11001000011010011110100110001100,
		32'b11001000000101101110100111000100,
		32'b11000111110000111110100111111101,
		32'b11000111011100001110101000110101,
		32'b11000111000111001110101001101101,
		32'b11000110110010011110101010100101,
		32'b11000110011101011110101011011100,
		32'b11000110001000011110101100010011,
		32'b11000101110011011110101101001010,
		32'b11000101011110001110101110000001,
		32'b11000101001001001110101110111000,
		32'b11000100110011111110101111101110,
		32'b11000100011110101110110000100100,
		32'b11000100001001011110110001011001,
		32'b11000011110100001110110010001111,
		32'b11000011011110111110110011000100,
		32'b11000011001001011110110011111001,
		32'b11000010110100001110110100101101,
		32'b11000010011110101110110101100010,
		32'b11000010001001001110110110010110,
		32'b11000001110011101110110111001010,
		32'b11000001011101111110110111111101,
		32'b11000001001000011110111000110000,
		32'b11000000110010101110111001100011,
		32'b11000000011100111110111010010110,
		32'b11000000000111011110111011001001,
		32'b10111111110001011110111011111011,
		32'b10111111011011101110111100101101,
		32'b10111111000101111110111101011111,
		32'b10111110101111111110111110010000,
		32'b10111110011010001110111111000001,
		32'b10111110000100001110111111110010,
		32'b10111101101110001111000000100011,
		32'b10111101011000001111000001010011,
		32'b10111101000001111111000010000011,
		32'b10111100101011111111000010110011,
		32'b10111100010101101111000011100010,
		32'b10111011111111011111000100010010,
		32'b10111011101001011111000101000001,
		32'b10111011010011001111000101101111,
		32'b10111010111100101111000110011110,
		32'b10111010100110011111000111001100,
		32'b10111010010000001111000111111010,
		32'b10111001111001101111001000100111,
		32'b10111001100011001111001001010101,
		32'b10111001001100101111001010000010,
		32'b10111000110110001111001010101111,
		32'b10111000011111101111001011011011,
		32'b10111000001001001111001100000111,
		32'b10110111110010101111001100110011,
		32'b10110111011011111111001101011111,
		32'b10110111000101001111001110001010,
		32'b10110110101110101111001110110101,
		32'b10110110010111111111001111100000,
		32'b10110110000001001111010000001011,
		32'b10110101101010001111010000110101,
		32'b10110101010011011111010001011111,
		32'b10110100111100101111010010001001,
		32'b10110100100101101111010010110010,
		32'b10110100001110101111010011011011,
		32'b10110011110111101111010100000100,
		32'b10110011100000101111010100101101,
		32'b10110011001001101111010101010101,
		32'b10110010110010101111010101111101,
		32'b10110010011011101111010110100101,
		32'b10110010000100011111010111001100,
		32'b10110001101101011111010111110100,
		32'b10110001010110001111011000011011,
		32'b10110000111110111111011001000001,
		32'b10110000100111101111011001101000,
		32'b10110000010000011111011010001110,
		32'b10101111111001001111011010110011,
		32'b10101111100001111111011011011001,
		32'b10101111001010011111011011111110,
		32'b10101110110011001111011100100011,
		32'b10101110011011101111011101000111,
		32'b10101110000100011111011101101100,
		32'b10101101101100111111011110010000,
		32'b10101101010101011111011110110100,
		32'b10101100111101111111011111010111,
		32'b10101100100110001111011111111010,
		32'b10101100001110101111100000011101,
		32'b10101011110111001111100001000000,
		32'b10101011011111011111100001100010,
		32'b10101011000111111111100010000100,
		32'b10101010110000001111100010100110,
		32'b10101010011000011111100011000111,
		32'b10101010000000101111100011101000,
		32'b10101001101000111111100100001001,
		32'b10101001010001001111100100101010,
		32'b10101000111001011111100101001010,
		32'b10101000100001101111100101101010,
		32'b10101000001001101111100110001010,
		32'b10100111110001111111100110101001,
		32'b10100111011001111111100111001000,
		32'b10100111000001111111100111100111,
		32'b10100110101010001111101000000101,
		32'b10100110010010001111101000100100,
		32'b10100101111010001111101001000010,
		32'b10100101100010001111101001011111,
		32'b10100101001010001111101001111101,
		32'b10100100110001111111101010011010,
		32'b10100100011001111111101010110110,
		32'b10100100000001111111101011010011,
		32'b10100011101001101111101011101111,
		32'b10100011010001011111101100001011,
		32'b10100010111001011111101100100110,
		32'b10100010100001001111101101000010,
		32'b10100010001000111111101101011101,
		32'b10100001110000101111101101110111,
		32'b10100001011000011111101110010010,
		32'b10100001000000001111101110101100,
		32'b10100000100111111111101111000101,
		32'b10100000001111101111101111011111,
		32'b10011111110111001111101111111000,
		32'b10011111011110111111110000010001,
		32'b10011111000110011111110000101001,
		32'b10011110101110001111110001000010,
		32'b10011110010101101111110001011010,
		32'b10011101111101011111110001110001,
		32'b10011101100100111111110010001001,
		32'b10011101001100011111110010100000,
		32'b10011100110011111111110010110111,
		32'b10011100011011011111110011001101,
		32'b10011100000010111111110011100011,
		32'b10011011101010011111110011111001,
		32'b10011011010001111111110100001111,
		32'b10011010111001001111110100100100,
		32'b10011010100000101111110100111001,
		32'b10011010001000001111110101001110,
		32'b10011001101111011111110101100010,
		32'b10011001010110111111110101110110,
		32'b10011000111110001111110110001010,
		32'b10011000100101101111110110011101,
		32'b10011000001100111111110110110000,
		32'b10010111110100001111110111000011,
		32'b10010111011011011111110111010110,
		32'b10010111000010101111110111101000,
		32'b10010110101010001111110111111010,
		32'b10010110010001011111111000001100,
		32'b10010101111000101111111000011101,
		32'b10010101011111111111111000101110,
		32'b10010101000110111111111000111111,
		32'b10010100101110001111111001001111,
		32'b10010100010101011111111001011111,
		32'b10010011111100101111111001101111,
		32'b10010011100011101111111001111111,
		32'b10010011001010111111111010001110,
		32'b10010010110010001111111010011101,
		32'b10010010011001001111111010101011,
		32'b10010010000000011111111010111010,
		32'b10010001100111011111111011001000,
		32'b10010001001110011111111011010101,
		32'b10010000110101101111111011100011,
		32'b10010000011100101111111011110000,
		32'b10010000000011101111111011111101,
		32'b10001111101010111111111100001001,
		32'b10001111010001111111111100010101,
		32'b10001110111000111111111100100001,
		32'b10001110011111111111111100101101,
		32'b10001110000110111111111100111000,
		32'b10001101101101111111111101000011,
		32'b10001101010100111111111101001101,
		32'b10001100111011111111111101011000,
		32'b10001100100010111111111101100010,
		32'b10001100001001111111111101101011,
		32'b10001011110000111111111101110101,
		32'b10001011010111111111111101111110,
		32'b10001010111110111111111110000111,
		32'b10001010100101111111111110001111,
		32'b10001010001100111111111110010111,
		32'b10001001110011101111111110011111,
		32'b10001001011010101111111110100111,
		32'b10001001000001101111111110101110,
		32'b10001000101000101111111110110101,
		32'b10001000001111011111111110111100,
		32'b10000111110110011111111111000010,
		32'b10000111011101011111111111001000,
		32'b10000111000100001111111111001110,
		32'b10000110101011001111111111010011,
		32'b10000110010001111111111111011000,
		32'b10000101111000111111111111011101,
		32'b10000101011111111111111111100001,
		32'b10000101000110101111111111100101,
		32'b10000100101101101111111111101001,
		32'b10000100010100011111111111101101,
		32'b10000011111011011111111111110000,
		32'b10000011100010001111111111110011,
		32'b10000011001001001111111111110110,
		32'b10000010101111111111111111111000,
		32'b10000010010110111111111111111010,
		32'b10000001111101101111111111111100,
		32'b10000001100100101111111111111101,
		32'b10000001001011011111111111111110,
		32'b10000000110010011111111111111111,
		32'b10000000011001001111111111111111,
		32'b10000000000000001111111111111111,
		32'b00000000011001001111111111111111,
		32'b00000000110010011111111111111111,
		32'b00000001001011011111111111111110,
		32'b00000001100100101111111111111101,
		32'b00000001111101101111111111111100,
		32'b00000010010110111111111111111010,
		32'b00000010101111111111111111111000,
		32'b00000011001001001111111111110110,
		32'b00000011100010001111111111110011,
		32'b00000011111011011111111111110000,
		32'b00000100010100011111111111101101,
		32'b00000100101101101111111111101001,
		32'b00000101000110101111111111100101,
		32'b00000101011111111111111111100001,
		32'b00000101111000111111111111011101,
		32'b00000110010001111111111111011000,
		32'b00000110101011001111111111010011,
		32'b00000111000100001111111111001110,
		32'b00000111011101011111111111001000,
		32'b00000111110110011111111111000010,
		32'b00001000001111011111111110111100,
		32'b00001000101000101111111110110101,
		32'b00001001000001101111111110101110,
		32'b00001001011010101111111110100111,
		32'b00001001110011101111111110011111,
		32'b00001010001100111111111110010111,
		32'b00001010100101111111111110001111,
		32'b00001010111110111111111110000111,
		32'b00001011010111111111111101111110,
		32'b00001011110000111111111101110101,
		32'b00001100001001111111111101101011,
		32'b00001100100010111111111101100010,
		32'b00001100111011111111111101011000,
		32'b00001101010100111111111101001101,
		32'b00001101101101111111111101000011,
		32'b00001110000110111111111100111000,
		32'b00001110011111111111111100101101,
		32'b00001110111000111111111100100001,
		32'b00001111010001111111111100010101,
		32'b00001111101010111111111100001001,
		32'b00010000000011101111111011111101,
		32'b00010000011100101111111011110000,
		32'b00010000110101101111111011100011,
		32'b00010001001110011111111011010101,
		32'b00010001100111011111111011001000,
		32'b00010010000000011111111010111010,
		32'b00010010011001001111111010101011,
		32'b00010010110010001111111010011101,
		32'b00010011001010111111111010001110,
		32'b00010011100011101111111001111111,
		32'b00010011111100101111111001101111,
		32'b00010100010101011111111001011111,
		32'b00010100101110001111111001001111,
		32'b00010101000110111111111000111111,
		32'b00010101011111111111111000101110,
		32'b00010101111000101111111000011101,
		32'b00010110010001011111111000001100,
		32'b00010110101010001111110111111010,
		32'b00010111000010101111110111101000,
		32'b00010111011011011111110111010110,
		32'b00010111110100001111110111000011,
		32'b00011000001100111111110110110000,
		32'b00011000100101101111110110011101,
		32'b00011000111110001111110110001010,
		32'b00011001010110111111110101110110,
		32'b00011001101111011111110101100010,
		32'b00011010001000001111110101001110,
		32'b00011010100000101111110100111001,
		32'b00011010111001001111110100100100,
		32'b00011011010001111111110100001111,
		32'b00011011101010011111110011111001,
		32'b00011100000010111111110011100011,
		32'b00011100011011011111110011001101,
		32'b00011100110011111111110010110111,
		32'b00011101001100011111110010100000,
		32'b00011101100100111111110010001001,
		32'b00011101111101011111110001110001,
		32'b00011110010101101111110001011010,
		32'b00011110101110001111110001000010,
		32'b00011111000110011111110000101001,
		32'b00011111011110111111110000010001,
		32'b00011111110111001111101111111000,
		32'b00100000001111101111101111011111,
		32'b00100000100111111111101111000101,
		32'b00100001000000001111101110101100,
		32'b00100001011000011111101110010010,
		32'b00100001110000101111101101110111,
		32'b00100010001000111111101101011101,
		32'b00100010100001001111101101000010,
		32'b00100010111001011111101100100110,
		32'b00100011010001011111101100001011,
		32'b00100011101001101111101011101111,
		32'b00100100000001111111101011010011,
		32'b00100100011001111111101010110110,
		32'b00100100110001111111101010011010,
		32'b00100101001010001111101001111101,
		32'b00100101100010001111101001011111,
		32'b00100101111010001111101001000010,
		32'b00100110010010001111101000100100,
		32'b00100110101010001111101000000101,
		32'b00100111000001111111100111100111,
		32'b00100111011001111111100111001000,
		32'b00100111110001111111100110101001,
		32'b00101000001001101111100110001010,
		32'b00101000100001101111100101101010,
		32'b00101000111001011111100101001010,
		32'b00101001010001001111100100101010,
		32'b00101001101000111111100100001001,
		32'b00101010000000101111100011101000,
		32'b00101010011000011111100011000111,
		32'b00101010110000001111100010100110,
		32'b00101011000111111111100010000100,
		32'b00101011011111011111100001100010,
		32'b00101011110111001111100001000000,
		32'b00101100001110101111100000011101,
		32'b00101100100110001111011111111010,
		32'b00101100111101111111011111010111,
		32'b00101101010101011111011110110100,
		32'b00101101101100111111011110010000,
		32'b00101110000100011111011101101100,
		32'b00101110011011101111011101000111,
		32'b00101110110011001111011100100011,
		32'b00101111001010011111011011111110,
		32'b00101111100001111111011011011001,
		32'b00101111111001001111011010110011,
		32'b00110000010000011111011010001110,
		32'b00110000100111101111011001101000,
		32'b00110000111110111111011001000001,
		32'b00110001010110001111011000011011,
		32'b00110001101101011111010111110100,
		32'b00110010000100011111010111001100,
		32'b00110010011011101111010110100101,
		32'b00110010110010101111010101111101,
		32'b00110011001001101111010101010101,
		32'b00110011100000101111010100101101,
		32'b00110011110111101111010100000100,
		32'b00110100001110101111010011011011,
		32'b00110100100101101111010010110010,
		32'b00110100111100101111010010001001,
		32'b00110101010011011111010001011111,
		32'b00110101101010001111010000110101,
		32'b00110110000001001111010000001011,
		32'b00110110010111111111001111100000,
		32'b00110110101110101111001110110101,
		32'b00110111000101001111001110001010,
		32'b00110111011011111111001101011111,
		32'b00110111110010101111001100110011,
		32'b00111000001001001111001100000111,
		32'b00111000011111101111001011011011,
		32'b00111000110110001111001010101111,
		32'b00111001001100101111001010000010,
		32'b00111001100011001111001001010101,
		32'b00111001111001101111001000100111,
		32'b00111010010000001111000111111010,
		32'b00111010100110011111000111001100,
		32'b00111010111100101111000110011110,
		32'b00111011010011001111000101101111,
		32'b00111011101001011111000101000001,
		32'b00111011111111011111000100010010,
		32'b00111100010101101111000011100010,
		32'b00111100101011111111000010110011,
		32'b00111101000001111111000010000011,
		32'b00111101011000001111000001010011,
		32'b00111101101110001111000000100011,
		32'b00111110000100001110111111110010,
		32'b00111110011010001110111111000001,
		32'b00111110101111111110111110010000,
		32'b00111111000101111110111101011111,
		32'b00111111011011101110111100101101,
		32'b00111111110001011110111011111011,
		32'b01000000000111011110111011001001,
		32'b01000000011100111110111010010110,
		32'b01000000110010101110111001100011,
		32'b01000001001000011110111000110000,
		32'b01000001011101111110110111111101,
		32'b01000001110011101110110111001010,
		32'b01000010001001001110110110010110,
		32'b01000010011110101110110101100010,
		32'b01000010110100001110110100101101,
		32'b01000011001001011110110011111001,
		32'b01000011011110111110110011000100,
		32'b01000011110100001110110010001111,
		32'b01000100001001011110110001011001,
		32'b01000100011110101110110000100100,
		32'b01000100110011111110101111101110,
		32'b01000101001001001110101110111000,
		32'b01000101011110001110101110000001,
		32'b01000101110011011110101101001010,
		32'b01000110001000011110101100010011,
		32'b01000110011101011110101011011100,
		32'b01000110110010011110101010100101,
		32'b01000111000111001110101001101101,
		32'b01000111011100001110101000110101,
		32'b01000111110000111110100111111101,
		32'b01001000000101101110100111000100,
		32'b01001000011010011110100110001100,
		32'b01001000101111001110100101010011,
		32'b01001001000011111110100100011001,
		32'b01001001011000011110100011100000,
		32'b01001001101101001110100010100110,
		32'b01001010000001101110100001101100,
		32'b01001010010110001110100000110010,
		32'b01001010101010011110011111110111,
		32'b01001010111110111110011110111101,
		32'b01001011010011001110011110000010,
		32'b01001011100111101110011101000110,
		32'b01001011111011111110011100001011,
		32'b01001100001111111110011011001111,
		32'b01001100100100001110011010010011,
		32'b01001100111000011110011001010111,
		32'b01001101001100011110011000011010,
		32'b01001101100000011110010111011101,
		32'b01001101110100011110010110100000,
		32'b01001110001000011110010101100011,
		32'b01001110011100001110010100100110,
		32'b01001110101111111110010011101000,
		32'b01001111000011111110010010101010,
		32'b01001111010111101110010001101100,
		32'b01001111101011001110010000101101,
		32'b01001111111110111110001111101111,
		32'b01010000010010011110001110110000,
		32'b01010000100101111110001101110001,
		32'b01010000111001011110001100110001,
		32'b01010001001100111110001011110010,
		32'b01010001100000011110001010110010,
		32'b01010001110011101110001001110001,
		32'b01010010000111001110001000110001,
		32'b01010010011010011110000111110001,
		32'b01010010101101011110000110110000,
		32'b01010011000000101110000101101111,
		32'b01010011010011101110000100101101,
		32'b01010011100110111110000011101100,
		32'b01010011111001111110000010101010,
		32'b01010100001100111110000001101000,
		32'b01010100011111101110000000100110,
		32'b01010100110010101101111111100011,
		32'b01010101000101011101111110100000,
		32'b01010101011000001101111101011110,
		32'b01010101101010111101111100011010,
		32'b01010101111101011101111011010111,
		32'b01010110010000001101111010010011,
		32'b01010110100010101101111001010000,
		32'b01010110110101001101111000001011,
		32'b01010111000111011101110111000111,
		32'b01010111011001111101110110000011,
		32'b01010111101100001101110100111110,
		32'b01010111111110011101110011111001,
		32'b01011000010000101101110010110100,
		32'b01011000100010111101110001101110,
		32'b01011000110101001101110000101001,
		32'b01011001000111001101101111100011,
		32'b01011001011001001101101110011101,
		32'b01011001101011001101101101010110,
		32'b01011001111100111101101100010000,
		32'b01011010001110111101101011001001,
		32'b01011010100000101101101010000010,
		32'b01011010110010011101101000111011,
		32'b01011011000100001101100111110011,
		32'b01011011010101101101100110101100,
		32'b01011011100111011101100101100100,
		32'b01011011111000111101100100011100,
		32'b01011100001010011101100011010100,
		32'b01011100011011101101100010001011,
		32'b01011100101101001101100001000010,
		32'b01011100111110011101011111111001,
		32'b01011101001111101101011110110000,
		32'b01011101100000111101011101100111,
		32'b01011101110001111101011100011101,
		32'b01011110000010111101011011010100,
		32'b01011110010100001101011010001010,
		32'b01011110100100111101011001000000,
		32'b01011110110101111101010111110101,
		32'b01011111000110101101010110101011,
		32'b01011111010111101101010101100000,
		32'b01011111101000001101010100010101,
		32'b01011111111000111101010011001010,
		32'b01100000001001101101010001111110,
		32'b01100000011010001101010000110011,
		32'b01100000101010101101001111100111,
		32'b01100000111011001101001110011011,
		32'b01100001001011011101001101001110,
		32'b01100001011011111101001100000010,
		32'b01100001101100001101001010110101,
		32'b01100001111100011101001001101001,
		32'b01100010001100011101001000011100,
		32'b01100010011100011101000111001110,
		32'b01100010101100101101000110000001,
		32'b01100010111100101101000100110011,
		32'b01100011001100011101000011100101,
		32'b01100011011100011101000010010111,
		32'b01100011101100001101000001001001,
		32'b01100011111011111100111111111011,
		32'b01100100001011011100111110101100,
		32'b01100100011011001100111101011110,
		32'b01100100101010101100111100001111,
		32'b01100100111010001100111010111111,
		32'b01100101001001101100111001110000,
		32'b01100101011000111100111000100001,
		32'b01100101101000001100110111010001,
		32'b01100101110111011100110110000001,
		32'b01100110000110101100110100110001,
		32'b01100110010101111100110011100001,
		32'b01100110100100111100110010010000,
		32'b01100110110011111100110000111111,
		32'b01100111000010111100101111101111,
		32'b01100111010001101100101110011110,
		32'b01100111100000101100101101001100,
		32'b01100111101111011100101011111011,
		32'b01100111111101111100101010101001,
		32'b01101000001100101100101001011000,
		32'b01101000011011001100101000000110,
		32'b01101000101001101100100110110100,
		32'b01101000111000001100100101100001,
		32'b01101001000110011100100100001111,
		32'b01101001010100111100100010111100,
		32'b01101001100011001100100001101001,
		32'b01101001110001001100100000010110,
		32'b01101001111111011100011111000011,
		32'b01101010001101011100011101110000,
		32'b01101010011011011100011100011100,
		32'b01101010101001011100011011001001,
		32'b01101010110111001100011001110101,
		32'b01101011000100111100011000100001,
		32'b01101011010010101100010111001101,
		32'b01101011100000011100010101111000,
		32'b01101011101110001100010100100100,
		32'b01101011111011101100010011001111,
		32'b01101100001001001100010001111010,
		32'b01101100010110011100010000100101,
		32'b01101100100011111100001111010000,
		32'b01101100110001001100001101111011,
		32'b01101100111110011100001100100101,
		32'b01101101001011011100001011010000,
		32'b01101101011000101100001001111010,
		32'b01101101100101101100001000100100,
		32'b01101101110010101100000111001110,
		32'b01101101111111011100000101110111,
		32'b01101110001100001100000100100001,
		32'b01101110011000111100000011001010,
		32'b01101110100101101100000001110011,
		32'b01101110110010011100000000011101,
		32'b01101110111110111011111111000101,
		32'b01101111001011011011111101101110,
		32'b01101111010111111011111100010111,
		32'b01101111100100001011111010111111,
		32'b01101111110000011011111001101000,
		32'b01101111111100101011111000010000,
		32'b01110000001000111011110110111000,
		32'b01110000010100111011110101100000,
		32'b01110000100000111011110100000111,
		32'b01110000101100111011110010101111,
		32'b01110000111000101011110001010110,
		32'b01110001000100101011101111111101,
		32'b01110001010000011011101110100101,
		32'b01110001011011111011101101001100,
		32'b01110001100111101011101011110010,
		32'b01110001110011001011101010011001,
		32'b01110001111110101011101001000000,
		32'b01110010001001111011100111100110,
		32'b01110010010101011011100110001100,
		32'b01110010100000101011100100110010,
		32'b01110010101011111011100011011000,
		32'b01110010110110111011100001111110,
		32'b01110011000001111011100000100100,
		32'b01110011001100111011011111001010,
		32'b01110011010111111011011101101111,
		32'b01110011100010101011011100010100,
		32'b01110011101101011011011010111010,
		32'b01110011111000001011011001011111,
		32'b01110100000010111011011000000100,
		32'b01110100001101011011010110101000,
		32'b01110100010111111011010101001101,
		32'b01110100100010011011010011110010,
		32'b01110100101100101011010010010110,
		32'b01110100110110111011010000111010,
		32'b01110101000001001011001111011110,
		32'b01110101001011011011001110000010,
		32'b01110101010101011011001100100110,
		32'b01110101011111011011001011001010,
		32'b01110101101001011011001001101110,
		32'b01110101110011001011001000010001,
		32'b01110101111101001011000110110101,
		32'b01110110000110111011000101011000,
		32'b01110110010000011011000011111011,
		32'b01110110011010001011000010011110,
		32'b01110110100011101011000001000001,
		32'b01110110101100111010111111100100,
		32'b01110110110110011010111110000111,
		32'b01110110111111101010111100101001,
		32'b01110111001000111010111011001100,
		32'b01110111010001111010111001101110,
		32'b01110111011011001010111000010001,
		32'b01110111100100001010110110110011,
		32'b01110111101101001010110101010101,
		32'b01110111110101111010110011110111,
		32'b01110111111110101010110010011000,
		32'b01111000000111011010110000111010,
		32'b01111000010000001010101111011100,
		32'b01111000011000101010101101111101,
		32'b01111000100001001010101100011111,
		32'b01111000101001101010101011000000,
		32'b01111000110001111010101001100001,
		32'b01111000111010001010101000000010,
		32'b01111001000010011010100110100011,
		32'b01111001001010101010100101000100,
		32'b01111001010010101010100011100101,
		32'b01111001011010101010100010000110,
		32'b01111001100010101010100000100110,
		32'b01111001101010011010011111000111,
		32'b01111001110010001010011101100111,
		32'b01111001111001111010011100000111,
		32'b01111010000001011010011010101000,
		32'b01111010001001001010011001001000,
		32'b01111010010000101010010111101000,
		32'b01111010010111111010010110001000,
		32'b01111010011111011010010100101000,
		32'b01111010100110101010010011000111,
		32'b01111010101101101010010001100111,
		32'b01111010110100111010010000000111,
		32'b01111010111011111010001110100110,
		32'b01111011000010111010001101000101,
		32'b01111011001001101010001011100101,
		32'b01111011010000101010001010000100,
		32'b01111011010111011010001000100011,
		32'b01111011011101111010000111000010,
		32'b01111011100100101010000101100001,
		32'b01111011101011001010000100000000,
		32'b01111011110001011010000010011111,
		32'b01111011110111111010000000111110,
		32'b01111011111110001001111111011100,
		32'b01111100000100011001111101111011,
		32'b01111100001010011001111100011001,
		32'b01111100010000101001111010111000,
		32'b01111100010110101001111001010110,
		32'b01111100011100011001110111110101,
		32'b01111100100010011001110110010011,
		32'b01111100101000001001110100110001,
		32'b01111100101101111001110011001111,
		32'b01111100110011011001110001101101,
		32'b01111100111000111001110000001011,
		32'b01111100111110011001101110101001,
		32'b01111101000011111001101101000111,
		32'b01111101001001001001101011100100,
		32'b01111101001110011001101010000010,
		32'b01111101010011101001101000100000,
		32'b01111101011000101001100110111101,
		32'b01111101011101101001100101011011,
		32'b01111101100010101001100011111000,
		32'b01111101100111011001100010010110,
		32'b01111101101100001001100000110011,
		32'b01111101110000111001011111010000,
		32'b01111101110101101001011101101101,
		32'b01111101111010001001011100001010,
		32'b01111101111110101001011010101000,
		32'b01111110000011001001011001000101,
		32'b01111110000111011001010111100010,
		32'b01111110001011101001010101111111,
		32'b01111110001111111001010100011011,
		32'b01111110010011111001010010111000,
		32'b01111110010111111001010001010101,
		32'b01111110011011111001001111110010,
		32'b01111110011111111001001110001110,
		32'b01111110100011101001001100101011,
		32'b01111110100111011001001011001000,
		32'b01111110101010111001001001100100,
		32'b01111110101110101001001000000001,
		32'b01111110110010001001000110011101,
		32'b01111110110101011001000100111001,
		32'b01111110111000111001000011010110,
		32'b01111110111100001001000001110010,
		32'b01111110111111011001000000001110,
		32'b01111111000010011000111110101011,
		32'b01111111000101011000111101000111,
		32'b01111111001000011000111011100011,
		32'b01111111001011011000111001111111,
		32'b01111111001110001000111000011011,
		32'b01111111010000111000110110110111,
		32'b01111111010011011000110101010011,
		32'b01111111010110001000110011101111,
		32'b01111111011000101000110010001011,
		32'b01111111011010111000110000100111,
		32'b01111111011101011000101111000011,
		32'b01111111011111101000101101011111,
		32'b01111111100001111000101011111011,
		32'b01111111100011111000101010010111,
		32'b01111111100101111000101000110011,
		32'b01111111100111111000100111001110,
		32'b01111111101001111000100101101010,
		32'b01111111101011101000100100000110,
		32'b01111111101101011000100010100010,
		32'b01111111101111001000100000111101,
		32'b01111111110000101000011111011001,
		32'b01111111110010001000011101110101,
		32'b01111111110011101000011100010000,
		32'b01111111110100111000011010101100,
		32'b01111111110110001000011001000111,
		32'b01111111110111011000010111100011,
		32'b01111111111000011000010101111111,
		32'b01111111111001011000010100011010,
		32'b01111111111010011000010010110110,
		32'b01111111111011011000010001010001,
		32'b01111111111100001000001111101101,
		32'b01111111111100111000001110001000,
		32'b01111111111101101000001100100100,
		32'b01111111111110001000001010111111,
		32'b01111111111110101000001001011011,
		32'b01111111111111001000000111110110,
		32'b01111111111111011000000110010010,
		32'b01111111111111101000000100101101,
		32'b01111111111111111000000011001001,
		32'b01111111111111111000000001100100};
				
		assign twiddle = ROM0[addr_t];

endmodule
